module tb_axi_slave_example;
	axi_slave_example

	AXI_LITE axi_lite ()
endmodule